/*
###############################################################################
# Copyright (c) 2019, PulseRain Technology LLC 
#
# This program is distributed under a dual license: an open source license, 
# and a commercial license. 
# 
# The open source license under which this program is distributed is the 
# GNU Public License version 3 (GPLv3).
#
# And for those who want to use this program in ways that are incompatible
# with the GPLv3, PulseRain Technology LLC offers commercial license instead.
# Please contact PulseRain Technology LLC (www.pulserain.com) for more detail.
#
###############################################################################
*/


//=============================================================================
// Remarks:
//     Top level wrapper for Onchip Debugger 
//=============================================================================

`include "debug_coprocessor.vh"

module debug_coprocessor_wrapper #(parameter BAUD_PERIOD=54) (
        input   wire                                clk,
        input   wire                                reset_n,
    
        
        input   wire                                RXD,
        output  wire                                TXD,
        
        input  wire                                                                 pram_read_enable_in,
        input  wire [`DEBUG_DATA_WIDTH * `DEBUG_FRAME_DATA_LEN - 1 : 0]             pram_read_data_in,
    
        output wire                                                                 pram_read_enable_out,
        output wire [`DEBUG_PRAM_ADDR_WIDTH - 3 : 0]                                pram_read_addr_out,
    
        
        output wire                                                                 pram_write_enable_out,
        output wire [`DEBUG_PRAM_ADDR_WIDTH - 3 : 0]                                pram_write_addr_out,
        output wire [`DEBUG_DATA_WIDTH * `DEBUG_FRAME_DATA_LEN  - 1 : 0]            pram_write_data_out,
        
        output wire                                                                 cpu_reset,
        output wire                                                                 cpu_start,
        output wire [`DEBUG_DATA_WIDTH * `DEBUG_FRAME_DATA_LEN - 1 : 0]             cpu_start_addr,
         
        output wire                                                                 debug_uart_tx_sel_ocd1_cpu0
    
);

    wire  [7 : 0]                                       SBUF_out;
    wire                                                TI, RI;
    
    wire                                                reply_enable;
    wire  [`DBG_NUM_OF_OPERATIONS - 1 : 0]              reply_debug_cmd;
    wire  [`DEBUG_ACK_PAYLOAD_BITS - 1 : 0]             reply_payload;
    
    wire                                                TX_done_pulse;
    
    wire                                                ctl_start_uart_tx;
    wire  [7 : 0]                                       SBUF_in;
    wire                                                reply_done;
    
    
   

    debug_UART #(.BAUD_PERIOD (BAUD_PERIOD)) debug_UART_i (
                .clk (clk),
                .reset_n (reset_n),
                .sync_reset (1'b0),
                .UART_enable (1'b1),
                .TX_enable_in (ctl_start_uart_tx),
                .RXD (RXD),
                .SBUF_in (SBUF_in),
                .REN (1'b1),
                .TXD (TXD),
                .SBUF_out (SBUF_out),
                .TX_done_pulse (TX_done_pulse), 
                .TI (TI),
                .RI (RI));
    
    debug_reply debug_reply_i (
            .clk (clk),
            .reset_n (reset_n),
            .reply_enable_in (reply_enable),
            .reply_debug_cmd (reply_debug_cmd),
            .reply_payload (reply_payload),
            
            .uart_tx_done (TX_done_pulse),
            
            .ctl_start_uart_tx (ctl_start_uart_tx),
            .uart_data_out (SBUF_in),
            .reply_done (reply_done));
    
    
    debug_coprocessor debug_coprocessor_i (
            .clk (clk),
            .reset_n (reset_n),
            .enable_in (RI),
            .debug_data_in (SBUF_out),
                        
            .reply_enable_out (reply_enable),
            .reply_debug_cmd (reply_debug_cmd),
            .reply_payload (reply_payload),
            
            .reply_done (reply_done),
            
            .pram_read_enable_in (pram_read_enable_in),
            .pram_read_data_in (pram_read_data_in),
            
            .pram_read_enable_out (pram_read_enable_out),
            .pram_read_addr_out (pram_read_addr_out),
            
            .pram_write_enable_out (pram_write_enable_out),
            .pram_write_addr_out (pram_write_addr_out),
            .pram_write_data_out (pram_write_data_out),
            
            .cpu_reset (cpu_reset),
            
            .cpu_start (cpu_start),
            .cpu_start_addr (cpu_start_addr),
    
            .debug_uart_tx_sel_ocd1_cpu0 (debug_uart_tx_sel_ocd1_cpu0)
    
            );
        
    
endmodule 

